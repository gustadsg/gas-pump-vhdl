-- teste --
Testando 123